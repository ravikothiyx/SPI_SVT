//////////////////////////////////////////////// 
// File:          spi_svt_inf.sv
// Version:       v1
// Developer:     Mayank
// Project Name:  SPI
// Discription:
/////////////////////////////////////////////////

interface spi_svt_inf();
endinterface : spi_svt_inf
