//////////////////////////////////////////////// 
// File:          spi_uvc_trans.sv
// Version:       v1
// Developer:     Harekrishna
// Project Name:  SPI
// Discription:
/////////////////////////////////////////////////


`ifndef SPI_UVC_TRANS_SV
`define SPI_UVC_TRANS_SV

class spi_uvc_trans extends uvm_sequence_item;
endclass
`endif 
