//////////////////////////////////////////////// 
// File:          spi_uvc_defines.sv
// Version:       v1
// Developer:     Mayank
// Project Name:  SPI
// Discription:
/////////////////////////////////////////////////


