//////////////////////////////////////////////// 
// File:          spi_uvc_inf.sv
// Version:       v1
// Developer:     Mayank
// Project Name:  SPI
// Discription:
/////////////////////////////////////////////////

interface spi_uvc_inf();
endinterface : spi_uvc_inf
