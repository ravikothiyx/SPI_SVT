//////////////////////////////////////////////// 
// File:          spi_svt_trans.sv
// Version:       v1
// Developer:     Harekrishna
// Project Name:  SPI
// Discription:
/////////////////////////////////////////////////


`ifndef SPI_SVT_TRANS_SV
`define SPI_SVT_TRANS_SV

class spi_svt_trans extends uvm_sequence_item;

endclass
`endif 
