//////////////////////////////////////////////// 
// File:          spi_uvc_defines.sv
// Version:       1.0
// Developer:     
// Project Name:  SPI
// Discription:
/////////////////////////////////////////////////


`define ADDR_WIDTH 8
`define DATA_WIDTH 8

