//////////////////////////////////////////////// 
// File:          spi_uvc_if.sv
// Version:       v1
// Developer:     Mayank
// Project Name:  SPI
// Discription:
/////////////////////////////////////////////////

interface spi_uvc_if();
endinterface : spi_uvc_if
