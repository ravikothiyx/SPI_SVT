///////////////////////////////////////////////
// File:          spi_uvc_seq_pkg.sv
// Version:       v1
// Developer:     Mayank
// Project Name:  SPI
// Discription:   SPI sequence package file 
/////////////////////////////////////////////////


/** Package Discription:*/


`ifndef SPI_UVC_SEQ_PKG_SV
`define SPI_UVC_SEQ_PKG_SV

package spi_uvc_seq_pkg;
   
   import uvm_pkg::*;
   `include "uvm_macros.svh"
   


endpackage : spi_uvc_seq_pkg
`endif /**SPI_UVC_SEQ_PKG*/
