///////////////////////////////////////////////
// File:          spi_uvc_master_pkg.sv
// Version:       v1
// Developer:     
// Project Name:  SPI
// Discription:   SPI master package file 
/////////////////////////////////////////////////


/** Package Discription:*/


`ifndef SPI_UVC_MASTER_PKG_SV
`define SPI_UVC_MASTER_PKG_SV

package spi_uvc_master_pkg;
   import uvm_pkg::*;
   `include "uvm_macros.svh"



endpackage : spi_uvc_master_pkg
`endif /**SPI_UVC_MASTER_PKG*/
