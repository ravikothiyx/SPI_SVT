//////////////////////////////////////////////// 
// File:          spi_svt_scoreboard.sv
// Version:       v1
// Developer:     Mayank
// Project Name:  SPI
// Discription:
/////////////////////////////////////////////////

`ifndef SPI_SVT_SCOREBOARD_SV
`define SPI_SVT_SCOREBOARD_SV

class spi_svt_scoreboard extends uvm_scoreboard;
   
   /** UVM Factory Registration Macro*/
   `uvm_component_utils(spi_svt_scoreboard);

   /** Transaction class instance*/
   spi_svt_trans trans_h;

   /** Analysis implementation for the master and slave monitor*/
   `uvm_analysis_imp_decl(_spi_svt_mstr_mon)
   `uvm_analysis_imp_decl(_spi_svt_slv_mon)

   /** Analysis implementation port declaration*/
   uvm_analysis_imp_spi_svt_mstr_mon#(spi_svt_trans,spi_svt_scoreboard) mstr_mon_imp;
   uvm_analysis_imp_spi_svt_slv_mon#(spi_svt_trans,spi_svt_scoreboard) slv_mon_imp;
   
   /** Standard UVM Methods*/
   extern function new(string name = "spi_svt_scoreboard",uvm_component parent);

   /** Write method of the master monitor*/
   extern function void write_spi_svt_mstr_mon(spi_svt_trans trans);

   /** Write method of the slave monitor*/
   extern function void write_spi_svt_slv_mon(spi_svt_trans trans);

   /** Run_phase*/
   extern task run_phase(uvm_phase phase);

endclass : spi_svt_scoreboard
`endif //: SPI_SVT_SCOREBOARD_SV

   /** Standard UVM Methods*/
   function spi_svt_scoreboard::new(string name = "spi_svt_scoreboard",uvm_component parent);
      super.new(name,parent);
     
      /** Constructing the implementation ports*/
      mstr_mon_imp = new("mstr_mon_imp",this);
      slv_mon_imp = new("slv_mon_imp",this);
   endfunction : new

   /** Write method of the master monitor*/
   function void spi_svt_scoreboard::write_spi_svt_mstr_mon(spi_svt_trans trans);
   endfunction : write_spi_svt_mstr_mon 

   /** Write method of the slave monitor*/
   function void spi_svt_scoreboard::write_spi_svt_slv_mon(spi_svt_trans trans);
   endfunction : write_spi_svt_slv_mon

   /** Run_phase*/
   task spi_svt_scoreboard::run_phase(uvm_phase phase);
      `uvm_info(get_type_name(),"START OF RUN_PHASE",UVM_HIGH);
      `uvm_info(get_type_name(),"INSIDE RUN_PHASE",UVM_DEBUG);
      `uvm_info(get_type_name(),"END OF RUN_PHASE",UVM_HIGH);
   endtask : run_phase
