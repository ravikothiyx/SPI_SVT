///////////////////////////////////////////////
// File:          spi_uvc_slave_pkg.sv
// Version:       v1
// Developer:     Mayank
// Project Name:  SPI
// Discription:   SPI slave package file 
/////////////////////////////////////////////////


/** Package Discription:*/


`ifndef SPI_UVC_PKG_SV
`define SPI_UVC_PKG_SV

package spi_uvc_slave_pkg;
    import uvm_pkg::*;
   `include "uvm_macros.svh"
  


 endpackage : spi_uvc_slave_pkg
`endif /**SPI_UVC_PKG*/
