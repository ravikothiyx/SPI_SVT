//////////////////////////////////////////////// 
// File:          spi_svt_top.sv
// Version:       v1
// Developer:     Mayank
// Project Name:  SPI
// Discription:
/////////////////////////////////////////////////


import uvm_pkg::*;
`include "uvm_macros.svh"

module spi_svt_top;
   

endmodule //spi_svt_top
